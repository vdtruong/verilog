`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:   13:50:11 04/23/2014 
// Design Name:   Van Truong
// Module Name:   GetPUCData 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 	This module collects data for the sdc host bus fifo.
//                         We need 1023 registers.  Whenever the host bus is
//                         ready for data, this module will increase to the next
//                         read address.
//									
//
//////////////////////////////////////////////////////////////////////////////////
module GetPUCData(
   input 					clk,
   input 					reset,	  
   output reg	[15:0]	rd_addr,			    // address to read data from bus arbitrator 
   output reg				rd_strb,			    // strobe to read data from bus arbitrator 
	// Data get packed into 64 bits word here.  Data from bus arbitrator. 
   input 		[35:0] 	rd_data,			    // data from bus arbitrator 
   input 					rd_rdy_strb,	    // strobe that data is ready	from b.a.  
   output reg	[63:0]	puc_data,		    // data for sdc fifo 
   output reg				puc_data_strb,		 // two clocks after rd_rdy_strb  
	input                rdy_for_nxt_pkt	 // ready for next packet (fifo_data) from puc.	  
   ); 
	 
	// Registers
	reg            rdy_for_nxt_pkt_z1;
	reg				rd_rdy_strb_z1;
	reg				rd_rdy_strb_z2;
	reg				puc_data_strb_z1;
	
	// Wires
	wire	[11:0]		sel_rd_addr;	// select which address to read
	
	// Initialize sequential logic
	initial			
	begin												
		rd_addr					   <= {16{1'b0}};			
		rd_strb					   <= 1'b0;
		puc_data					   <= {64{1'b0}};
		rdy_for_nxt_pkt_z1    	<= 1'b0;
		rd_rdy_strb_z1		 	   <= 1'b0;
		rd_rdy_strb_z2		 	   <= 1'b0;
		puc_data_strb			 	<= 1'b0;
		puc_data_strb_z1		 	<= 1'b0;
	end     
	
	// Create delays.
	always@(posedge clk)
	begin
		if (reset) begin
		   rdy_for_nxt_pkt_z1    	<= 1'b0;
			rd_rdy_strb_z1		 	   <= 1'b0;
			rd_rdy_strb_z2		 	   <= 1'b0;
			puc_data_strb			 	<= 1'b0;
			puc_data_strb_z1		 	<= 1'b0;
		end
		else begin  
		   rdy_for_nxt_pkt_z1    	<= rdy_for_nxt_pkt;
			rd_rdy_strb_z1		 	   <= rd_rdy_strb;
			rd_rdy_strb_z2		 	   <= rd_rdy_strb_z1;
			puc_data_strb			 	<= rd_rdy_strb_z2;
			puc_data_strb_z1		 	<= puc_data_strb;
		end
	end
  
	//---------------------------------------------------------------
	// Counts to 1024 addresses.
	//
	defparam ADDR_COUNTER.dw 	= 12;
	defparam ADDR_COUNTER.max 	= 12'h400; 
	//---------------------------------------------------------------
	Counter ADDR_COUNTER 
	(
		.clk(clk),
		.reset(reset),
		// Get a new address
		// every time we send away the packet to
		// the fifo.
		.enable(rdy_for_nxt_pkt),
		.cntr(sel_rd_addr),
		.strb()
	);		
	
	// Strobe to read after we have increased the address.
	always@(posedge clk)
	begin
		if (reset) 
			rd_strb 	<= 1'b0;
		else if (rdy_for_nxt_pkt_z1) 	// may need to delay more     
			rd_strb 	<= 1'b1;				// read from bus arbitrator
		else  
			rd_strb 	<= 1'b0;
	end
	
	always@(posedge clk)
	begin
		if (reset) 
			puc_data		<= {64{1'b0}};
		else if (rd_rdy_strb)     
			puc_data		<= {{28{1'b0}},rd_data};
		else  
			puc_data		<= puc_data;
	end
	
	// Select which address to read base on counter.
   always @(sel_rd_addr)
      case (sel_rd_addr)
         12'h001: 	rd_addr = 16'h0000;
         12'h002: 	rd_addr = 16'h0001;
         12'h003: 	rd_addr = 16'h0002;
         12'h004: 	rd_addr = 16'h0003;
         12'h005: 	rd_addr = 16'h0004;
         12'h006: 	rd_addr = 16'h0005;
         12'h007: 	rd_addr = 16'h0006;
         12'h008: 	rd_addr = 16'h0007;
         12'h009: 	rd_addr = 16'h0008;
         12'h00A: 	rd_addr = 16'h0009;
         12'h00B: 	rd_addr = 16'h000A;
         12'h00C: 	rd_addr = 16'h000B;
         12'h00D: 	rd_addr = 16'h000C;
         12'h00E: 	rd_addr = 16'h000D;
         12'h00F: 	rd_addr = 16'h000E;
         12'h010: 	rd_addr = 16'h000F;
         12'h011: 	rd_addr = 16'h0010;
         12'h012: 	rd_addr = 16'h0011;
         12'h013: 	rd_addr = 16'h0012;
         12'h014: 	rd_addr = 16'h0013;
         12'h015: 	rd_addr = 16'h0014;
         12'h016: 	rd_addr = 16'h0015;
         12'h017: 	rd_addr = 16'h0016;
         12'h018: 	rd_addr = 16'h0017;
         12'h019: 	rd_addr = 16'h0018;
         12'h01A: 	rd_addr = 16'h0019;
         12'h01B: 	rd_addr = 16'h001A;
         12'h01C: 	rd_addr = 16'h001B;
         12'h01D: 	rd_addr = 16'h001C;
         12'h01E: 	rd_addr = 16'h001D;
         12'h01F: 	rd_addr = 16'h001E;
         12'h020: 	rd_addr = 16'h001F;
         12'h021: 	rd_addr = 16'h0020;
         12'h022: 	rd_addr = 16'h0021;
         12'h023: 	rd_addr = 16'h0022;
         12'h024: 	rd_addr = 16'h0023;
         12'h025: 	rd_addr = 16'h0024;
         12'h026: 	rd_addr = 16'h0025;
         12'h027: 	rd_addr = 16'h0026;
         12'h028: 	rd_addr = 16'h0027;
         12'h029: 	rd_addr = 16'h0028;
         12'h02A: 	rd_addr = 16'h0029;
         12'h02B: 	rd_addr = 16'h002A;
         12'h02C: 	rd_addr = 16'h002B;
         12'h02D: 	rd_addr = 16'h002C;
         12'h02E: 	rd_addr = 16'h002D;
         12'h02F: 	rd_addr = 16'h002E;
         12'h030: 	rd_addr = 16'h002F;
         12'h031: 	rd_addr = 16'h0030;
         12'h032: 	rd_addr = 16'h0031;
         12'h033: 	rd_addr = 16'h0032;
         12'h034: 	rd_addr = 16'h0033;
         12'h035: 	rd_addr = 16'h0034;
         12'h036: 	rd_addr = 16'h0035;
         12'h037: 	rd_addr = 16'h0036;
         12'h038: 	rd_addr = 16'h0037;
         12'h039: 	rd_addr = 16'h0038;
         12'h03A: 	rd_addr = 16'h0039;
         12'h03B: 	rd_addr = 16'h003A;
         12'h03C: 	rd_addr = 16'h003B;
         12'h03D: 	rd_addr = 16'h003C;
         12'h03E: 	rd_addr = 16'h003D;
         12'h03F: 	rd_addr = 16'h003E;
         12'h040: 	rd_addr = 16'h003F;
         12'h041: 	rd_addr = 16'h0040;
         12'h042: 	rd_addr = 16'h0041;
         12'h043: 	rd_addr = 16'h0042;
         12'h044: 	rd_addr = 16'h0043;
         12'h045: 	rd_addr = 16'h0044;
         12'h046: 	rd_addr = 16'h0045;
         12'h047: 	rd_addr = 16'h0046;
         12'h048: 	rd_addr = 16'h0047;
         12'h049: 	rd_addr = 16'h0048;
         12'h04A: 	rd_addr = 16'h0049;
         12'h04B: 	rd_addr = 16'h004A;
         12'h04C: 	rd_addr = 16'h004B;
         12'h04D: 	rd_addr = 16'h004C;
         12'h04E: 	rd_addr = 16'h004D;
         12'h04F: 	rd_addr = 16'h004E;
         12'h050: 	rd_addr = 16'h004F;
         12'h051: 	rd_addr = 16'h0050;
         12'h052: 	rd_addr = 16'h0051;
         12'h053: 	rd_addr = 16'h0052;
         12'h054: 	rd_addr = 16'h0053;
         12'h055: 	rd_addr = 16'h0054;
         12'h056: 	rd_addr = 16'h0055;
         12'h057: 	rd_addr = 16'h0056;
         12'h058: 	rd_addr = 16'h0057;
         12'h059: 	rd_addr = 16'h0058;
         12'h05A: 	rd_addr = 16'h0059;
         12'h05B: 	rd_addr = 16'h005A;
         12'h05C: 	rd_addr = 16'h005B;
         12'h05D: 	rd_addr = 16'h005C;
         12'h05E: 	rd_addr = 16'h005D;
         12'h05F: 	rd_addr = 16'h005E;
         12'h060: 	rd_addr = 16'h005F;
         12'h061: 	rd_addr = 16'h0060;
         12'h062: 	rd_addr = 16'h0061;
         12'h063: 	rd_addr = 16'h0062;
         12'h064:    rd_addr = 16'h0063;
         12'h065:    rd_addr = 16'h0064;
         12'h066:    rd_addr = 16'h0065;
         12'h067:    rd_addr = 16'h0066; 	
         12'h068:    rd_addr = 16'h0067;	
         12'h069:    rd_addr = 16'h0068;	
         12'h06A: 	rd_addr = 16'h0069;
         12'h06B: 	rd_addr = 16'h006A;
         12'h06C: 	rd_addr = 16'h006B;
         12'h06D: 	rd_addr = 16'h006C;
         12'h06E: 	rd_addr = 16'h006D;
         12'h06F: 	rd_addr = 16'h006E;
         12'h070:    rd_addr = 16'h006F;
         12'h071: 	rd_addr = 16'h0070;
         12'h072: 	rd_addr = 16'h0071;
         12'h073: 	rd_addr = 16'h0072;
         12'h074: 	rd_addr = 16'h0073;
         12'h075: 	rd_addr = 16'h0074;
         12'h076:    rd_addr = 16'h0075;
         12'h077:    rd_addr = 16'h0076; 	
         12'h078:    rd_addr = 16'h0077;	
         12'h079:    rd_addr = 16'h0078;	
         12'h07A:    rd_addr = 16'h0079;	
         12'h07B:    rd_addr = 16'h007A;	
         12'h07C:    rd_addr = 16'h007B;	
         12'h07D: 	rd_addr = 16'h007C;
         12'h07E: 	rd_addr = 16'h007D;
         12'h07F: 	rd_addr = 16'h007E;
         12'h080:    rd_addr = 16'h007F;
         12'h081: 	rd_addr = 16'h0080;
         12'h082: 	rd_addr = 16'h0081;
         12'h083: 	rd_addr = 16'h0082;
         12'h084: 	rd_addr = 16'h0083;
         12'h085: 	rd_addr = 16'h0084;
         12'h086:    rd_addr = 16'h0085;
         12'h087:  	rd_addr = 16'h0086;
         12'h088: 	rd_addr = 16'h0087;
         12'h089: 	rd_addr = 16'h0088;
         12'h08A: 	rd_addr = 16'h0089;
         12'h08B: 	rd_addr = 16'h008A;
         12'h08C: 	rd_addr = 16'h008B;
         12'h08D: 	rd_addr = 16'h008C;
         12'h08E:    rd_addr = 16'h008D;	
         12'h08F: 	rd_addr = 16'h008E;
         12'h090:    rd_addr = 16'h008F;
         12'h091: 	rd_addr = 16'h0090;
         12'h092: 	rd_addr = 16'h0091;
         12'h093: 	rd_addr = 16'h0092;
         12'h094: 	rd_addr = 16'h0093;
         12'h095: 	rd_addr = 16'h0094;
         12'h096:    rd_addr = 16'h0095;
         12'h097:    rd_addr = 16'h0096;  	
         12'h098: 	rd_addr = 16'h0097;
         12'h099: 	rd_addr = 16'h0098;
         12'h09A: 	rd_addr = 16'h0099;
         12'h09B:    rd_addr = 16'h009A;	
         12'h09C:    rd_addr = 16'h009B; 	
         12'h09D: 	rd_addr = 16'h009C;
         12'h09E: 	rd_addr = 16'h009D;
         12'h09F: 	rd_addr = 16'h009E;
         12'h0A0:    rd_addr = 16'h009F;
         12'h0A1: 	rd_addr = 16'h00A0;
         12'h0A2: 	rd_addr = 16'h00A1;
         12'h0A3: 	rd_addr = 16'h00A2;
         12'h0A4:    rd_addr = 16'h00A3;	
         12'h0A5:    rd_addr = 16'h00A4;	
         12'h0A6:    rd_addr = 16'h00A5;
         12'h0A7:  	rd_addr = 16'h00A6;
         12'h0A8: 	rd_addr = 16'h00A7;
         12'h0A9: 	rd_addr = 16'h00A8;
         12'h0AA: 	rd_addr = 16'h00A9;
         12'h0AB: 	rd_addr = 16'h00AA;
         12'h0AC: 	rd_addr = 16'h00AB;
         12'h0AD: 	rd_addr = 16'h00AC;
         12'h0AE: 	rd_addr = 16'h00AD;
         12'h0AF: 	rd_addr = 16'h00AE;
         12'h0B0: 	rd_addr = 16'h00AF;
         12'h0B1: 	rd_addr = 16'h00B0;
         12'h0B2: 	rd_addr = 16'h00B1;
         12'h0B3: 	rd_addr = 16'h00B2;
         12'h0B4: 	rd_addr = 16'h00B3;
         12'h0B5:    rd_addr = 16'h00B4;
         12'h0B6:  	rd_addr = 16'h00B5;
         12'h0B7:    rd_addr = 16'h00B6;	
         12'h0B8: 	rd_addr = 16'h00B7;
         12'h0B9: 	rd_addr = 16'h00B8;
         12'h0BA: 	rd_addr = 16'h00B9;
         12'h0BB:    rd_addr = 16'h00BA;   	
         12'h0BC:    rd_addr = 16'h00BB;
         12'h0BD:    rd_addr = 16'h00BC;	
         12'h0BE: 	rd_addr = 16'h00BD;
         12'h0BF: 	rd_addr = 16'h00BE;
         12'h0C0: 	rd_addr = 16'h00BF;
         12'h0C1: 	rd_addr = 16'h00C0;
         12'h0C2: 	rd_addr = 16'h00C1;
         12'h0C3: 	rd_addr = 16'h00C2;
         12'h0C4: 	rd_addr = 16'h00C3;
         12'h0C5:    rd_addr = 16'h00C4;
         12'h0C6:  	rd_addr = 16'h00C5;
         12'h0C7: 	rd_addr = 16'h00C6;
         12'h0C8: 	rd_addr = 16'h00C7;
         12'h0C9: 	rd_addr = 16'h00C8;
         12'h0CA: 	rd_addr = 16'h00C9;
         12'h0CB: 	rd_addr = 16'h00CA;
         12'h0CC: 	rd_addr = 16'h00CB;
         12'h0CD:    rd_addr = 16'h00CC;	
         12'h0CE:    rd_addr = 16'h00CD;	
         12'h0CF: 	rd_addr = 16'h00CE;
         12'h0D0:    rd_addr = 16'h00CF;	
         12'h0D1: 	rd_addr = 16'h00D0;
         12'h0D2: 	rd_addr = 16'h00D1;
         12'h0D3: 	rd_addr = 16'h00D2;
         12'h0D4: 	rd_addr = 16'h00D3;
         12'h0D5:    rd_addr = 16'h00D4;
         12'h0D6:  	rd_addr = 16'h00D5;
         12'h0D7: 	rd_addr = 16'h00D6;
         12'h0D8: 	rd_addr = 16'h00D7;
         12'h0D9: 	rd_addr = 16'h00D8;
         12'h0DA: 	rd_addr = 16'h00D9;
         12'h0DB: 	rd_addr = 16'h00DA;
         12'h0DC: 	rd_addr = 16'h00DB;
         12'h0DD: 	rd_addr = 16'h00DC;
         12'h0DE: 	rd_addr = 16'h00DD;
         12'h0DF: 	rd_addr = 16'h00DE;
         12'h0E0: 	rd_addr = 16'h00DF;
         12'h0E1: 	rd_addr = 16'h00E0;
         12'h0E2: 	rd_addr = 16'h00E1;
         12'h0E3:    rd_addr = 16'h00E2;	
         12'h0E4: 	rd_addr = 16'h00E3;
         12'h0E5:    rd_addr = 16'h00E4; 
         12'h0E6:  	rd_addr = 16'h00E5;
         12'h0E7: 	rd_addr = 16'h00E6;
         12'h0E8: 	rd_addr = 16'h00E7;
         12'h0E9: 	rd_addr = 16'h00E8;
         12'h0EA: 	rd_addr = 16'h00E9;
         12'h0EB: 	rd_addr = 16'h00EA;
         12'h0EC: 	rd_addr = 16'h00EB;
         12'h0ED: 	rd_addr = 16'h00EC;
         12'h0EE: 	rd_addr = 16'h00ED;
         12'h0EF: 	rd_addr = 16'h00EE;
         12'h0F0: 	rd_addr = 16'h00EF;
         12'h0F1: 	rd_addr = 16'h00F0;
         12'h0F2: 	rd_addr = 16'h00F1;
         12'h0F3: 	rd_addr = 16'h00F2;
         12'h0F4: 	rd_addr = 16'h00F3;
         12'h0F5:    rd_addr = 16'h00F4;
         12'h0F6:  	rd_addr = 16'h00F5;
         12'h0F7: 	rd_addr = 16'h00F6;
         12'h0F8: 	rd_addr = 16'h00F7;
         12'h0F9: 	rd_addr = 16'h00F8;
         12'h0FA: 	rd_addr = 16'h00F9;
         12'h0FB: 	rd_addr = 16'h00FA;
         12'h0FC: 	rd_addr = 16'h00FB;
         12'h0FD: 	rd_addr = 16'h00FC;
         12'h0FE: 	rd_addr = 16'h00FD;
         12'h0FF: 	rd_addr = 16'h00FE;
         12'h100:    rd_addr = 16'h00FF;
         12'h101: 	rd_addr = 16'h0100;
         12'h102: 	rd_addr = 16'h0101;
         12'h103: 	rd_addr = 16'h0102;
         12'h104: 	rd_addr = 16'h0103;
         12'h105: 	rd_addr = 16'h0104;
         12'h106: 	rd_addr = 16'h0105;
         12'h107: 	rd_addr = 16'h0106;
         12'h108: 	rd_addr = 16'h0107;
         12'h109: 	rd_addr = 16'h0108;
         12'h10A: 	rd_addr = 16'h0109;
         12'h10B: 	rd_addr = 16'h010A;
         12'h10C: 	rd_addr = 16'h010B;
         12'h10D: 	rd_addr = 16'h010C;
         12'h10E: 	rd_addr = 16'h010D;
         12'h10F: 	rd_addr = 16'h010E;
         12'h110: 	rd_addr = 16'h010F;
         12'h111: 	rd_addr = 16'h0110;
         12'h112: 	rd_addr = 16'h0111;
         12'h113: 	rd_addr = 16'h0112;
         12'h114: 	rd_addr = 16'h0113;
         12'h115: 	rd_addr = 16'h0114;
         12'h116: 	rd_addr = 16'h0115;
         12'h117: 	rd_addr = 16'h0116;
         12'h118: 	rd_addr = 16'h0117;
         12'h119: 	rd_addr = 16'h0118;
         12'h11A: 	rd_addr = 16'h0119;
         12'h11B: 	rd_addr = 16'h011A;
         12'h11C: 	rd_addr = 16'h011B;
         12'h11D: 	rd_addr = 16'h011C;
         12'h11E: 	rd_addr = 16'h011D;
         12'h11F: 	rd_addr = 16'h011E;
         12'h120: 	rd_addr = 16'h011F;
         12'h121: 	rd_addr = 16'h0120;
         12'h122: 	rd_addr = 16'h0121;
         12'h123: 	rd_addr = 16'h0122;
         12'h124: 	rd_addr = 16'h0123;
         12'h125: 	rd_addr = 16'h0124;
         12'h126: 	rd_addr = 16'h0125;
         12'h127: 	rd_addr = 16'h0126;
         12'h128: 	rd_addr = 16'h0127;
         12'h129: 	rd_addr = 16'h0128;
         12'h12A: 	rd_addr = 16'h0129;
         12'h12B: 	rd_addr = 16'h012A;
         12'h12C: 	rd_addr = 16'h012B;
         12'h12D: 	rd_addr = 16'h012C;
         12'h12E: 	rd_addr = 16'h012D;
         12'h12F: 	rd_addr = 16'h012E;
         12'h130: 	rd_addr = 16'h012F;
         12'h131: 	rd_addr = 16'h0130;
         12'h132: 	rd_addr = 16'h0131;
         12'h133: 	rd_addr = 16'h0132;
         12'h134: 	rd_addr = 16'h0133;
         12'h135: 	rd_addr = 16'h0134;
         12'h136: 	rd_addr = 16'h0135;
         12'h137: 	rd_addr = 16'h0136;
         12'h138: 	rd_addr = 16'h0137;
         12'h139: 	rd_addr = 16'h0138;
         12'h13A: 	rd_addr = 16'h0139;
         12'h13B: 	rd_addr = 16'h013A;
         12'h13C: 	rd_addr = 16'h013B;
         12'h13D: 	rd_addr = 16'h013C;
         12'h13E: 	rd_addr = 16'h013D;
         12'h13F: 	rd_addr = 16'h013E;
         12'h140: 	rd_addr = 16'h013F;
         12'h141: 	rd_addr = 16'h0140;
         12'h142: 	rd_addr = 16'h0141;
         12'h143: 	rd_addr = 16'h0142;
         12'h144: 	rd_addr = 16'h0143;
         12'h145: 	rd_addr = 16'h0144;
         12'h146: 	rd_addr = 16'h0145;
         12'h147: 	rd_addr = 16'h0146;
         12'h148: 	rd_addr = 16'h0147;
         12'h149: 	rd_addr = 16'h0148;
         12'h14A: 	rd_addr = 16'h0149;
         12'h14B: 	rd_addr = 16'h014A;
         12'h14C: 	rd_addr = 16'h014B;
         12'h14D: 	rd_addr = 16'h014C;
         12'h14E: 	rd_addr = 16'h014D;
         12'h14F: 	rd_addr = 16'h014E;
         12'h150: 	rd_addr = 16'h014F;
         12'h151: 	rd_addr = 16'h0150;
         12'h152: 	rd_addr = 16'h0151;
         12'h153: 	rd_addr = 16'h0152;
         12'h154: 	rd_addr = 16'h0153;
         12'h155: 	rd_addr = 16'h0154;
         12'h156: 	rd_addr = 16'h0155;
         12'h157: 	rd_addr = 16'h0156;
         12'h158: 	rd_addr = 16'h0157;
         12'h159: 	rd_addr = 16'h0158;
         12'h15A: 	rd_addr = 16'h0159;
         12'h15B: 	rd_addr = 16'h015A;
         12'h15C: 	rd_addr = 16'h015B;
         12'h15D: 	rd_addr = 16'h015C;
         12'h15E: 	rd_addr = 16'h015D;
         12'h15F: 	rd_addr = 16'h015E;
         12'h160: 	rd_addr = 16'h015F;
         12'h161: 	rd_addr = 16'h0160;
         12'h162: 	rd_addr = 16'h0161;
         12'h163:    rd_addr = 16'h0162;    
         12'h164:    rd_addr = 16'h0163;    
         12'h165:    rd_addr = 16'h0164;    
         12'h166:    rd_addr = 16'h0165;    
         12'h167:  	rd_addr = 16'h0166;    
         12'h168: 	rd_addr = 16'h0167;      
         12'h169: 	rd_addr = 16'h0168;      
         12'h16A: 	rd_addr = 16'h0169;      
         12'h16B: 	rd_addr = 16'h016A;      
         12'h16C: 	rd_addr = 16'h016B;      
         12'h16D: 	rd_addr = 16'h016C;      
         12'h16E: 	rd_addr = 16'h016D;      
         12'h16F: 	rd_addr = 16'h016E;      
         12'h170:    rd_addr = 16'h016F;      
         12'h171: 	rd_addr = 16'h0170;      
         12'h172: 	rd_addr = 16'h0171;      
         12'h173: 	rd_addr = 16'h0172;      
         12'h174: 	rd_addr = 16'h0173;      
         12'h175: 	rd_addr = 16'h0174;      
         12'h176:    rd_addr = 16'h0175;      
         12'h177:  	rd_addr = 16'h0176;      
         12'h178: 	rd_addr = 16'h0177;      
         12'h179: 	rd_addr = 16'h0178;
         12'h17A:    rd_addr = 16'h0179;         	
         12'h17B:    rd_addr = 16'h017A;      	
         12'h17C: 	rd_addr = 16'h017B;
         12'h17D: 	rd_addr = 16'h017C;
         12'h17E: 	rd_addr = 16'h017D;
         12'h17F: 	rd_addr = 16'h017E;
         12'h180:    rd_addr = 16'h017F;
         12'h181: 	rd_addr = 16'h0180;
         12'h182: 	rd_addr = 16'h0181;
         12'h183: 	rd_addr = 16'h0182;
         12'h184: 	rd_addr = 16'h0183;
         12'h185: 	rd_addr = 16'h0184;
         12'h186:    rd_addr = 16'h0185;
         12'h187:  	rd_addr = 16'h0186;
         12'h188: 	rd_addr = 16'h0187;
         12'h189: 	rd_addr = 16'h0188;
         12'h18A: 	rd_addr = 16'h0189;
         12'h18B: 	rd_addr = 16'h018A;
         12'h18C: 	rd_addr = 16'h018B;
         12'h18D: 	rd_addr = 16'h018C;
         12'h18E: 	rd_addr = 16'h018D;
         12'h18F: 	rd_addr = 16'h018E;
         12'h190:    rd_addr = 16'h018F;   
         12'h191:    rd_addr = 16'h0190;   	
         12'h192: 	rd_addr = 16'h0191;
         12'h193: 	rd_addr = 16'h0192;
         12'h194: 	rd_addr = 16'h0193;
         12'h195: 	rd_addr = 16'h0194;
         12'h196:    rd_addr = 16'h0195;
         12'h197:  	rd_addr = 16'h0196;
         12'h198: 	rd_addr = 16'h0197;
         12'h199: 	rd_addr = 16'h0198;
         12'h19A: 	rd_addr = 16'h0199;
         12'h19B:    rd_addr = 16'h019A;	      
         12'h19C: 	rd_addr = 16'h019B;      
         12'h19D: 	rd_addr = 16'h019C;      
         12'h19E: 	rd_addr = 16'h019D;      
         12'h19F: 	rd_addr = 16'h019E;      
         12'h1A0:    rd_addr = 16'h019F;      
         12'h1A1:    rd_addr = 16'h01A0;            	
         12'h1A2:    rd_addr = 16'h01A1;   	
         12'h1A3: 	rd_addr = 16'h01A2;      
         12'h1A4: 	rd_addr = 16'h01A3;      
         12'h1A5: 	rd_addr = 16'h01A4;      
         12'h1A6:    rd_addr = 16'h01A5;      
         12'h1A7:  	rd_addr = 16'h01A6;      
         12'h1A8: 	rd_addr = 16'h01A7;      
         12'h1A9: 	rd_addr = 16'h01A8;      
         12'h1AA: 	rd_addr = 16'h01A9;      
         12'h1AB: 	rd_addr = 16'h01AA;      
         12'h1AC: 	rd_addr = 16'h01AB;      
         12'h1AD: 	rd_addr = 16'h01AC;      
         12'h1AE: 	rd_addr = 16'h01AD;      
         12'h1AF: 	rd_addr = 16'h01AE;      
         12'h1B0: 	rd_addr = 16'h01AF;      
         12'h1B1: 	rd_addr = 16'h01B0;      
         12'h1B2: 	rd_addr = 16'h01B1;      
         12'h1B3: 	rd_addr = 16'h01B2;      
         12'h1B4: 	rd_addr = 16'h01B3;      
         12'h1B5:    rd_addr = 16'h01B4;      
         12'h1B6:  	rd_addr = 16'h01B5;      
         12'h1B7: 	rd_addr = 16'h01B6;      
         12'h1B8: 	rd_addr = 16'h01B7;      
         12'h1B9: 	rd_addr = 16'h01B8;      
         12'h1BA: 	rd_addr = 16'h01B9;      
         12'h1BB:    rd_addr = 16'h01BA;      	
         12'h1BC:  	rd_addr = 16'h01BB;      
         12'h1BD: 	rd_addr = 16'h01BC;      
         12'h1BE: 	rd_addr = 16'h01BD;      
         12'h1BF: 	rd_addr = 16'h01BE;      
         12'h1C0: 	rd_addr = 16'h01BF;      
         12'h1C1: 	rd_addr = 16'h01C0;      
         12'h1C2: 	rd_addr = 16'h01C1;      
         12'h1C3: 	rd_addr = 16'h01C2;      
         12'h1C4: 	rd_addr = 16'h01C3;      
         12'h1C5:    rd_addr = 16'h01C4;      
         12'h1C6:    rd_addr = 16'h01C5;      
         12'h1C7: 	rd_addr = 16'h01C6;      
         12'h1C8: 	rd_addr = 16'h01C7;      
         12'h1C9: 	rd_addr = 16'h01C8;      
         12'h1CA: 	rd_addr = 16'h01C9;      
         12'h1CB: 	rd_addr = 16'h01CA;      
         12'h1CC: 	rd_addr = 16'h01CB;      
         12'h1CD: 	rd_addr = 16'h01CC;      
         12'h1CE: 	rd_addr = 16'h01CD;      
         12'h1CF: 	rd_addr = 16'h01CE;      
         12'h1D0: 	rd_addr = 16'h01CF;      
         12'h1D1: 	rd_addr = 16'h01D0;      
         12'h1D2: 	rd_addr = 16'h01D1;      
         12'h1D3: 	rd_addr = 16'h01D2;      
         12'h1D4: 	rd_addr = 16'h01D3;      
         12'h1D5:    rd_addr = 16'h01D4;      
         12'h1D6:    rd_addr = 16'h01D5;      
         12'h1D7:    rd_addr = 16'h01D6;      	
         12'h1D8: 	rd_addr = 16'h01D7;      
         12'h1D9: 	rd_addr = 16'h01D8;      
         12'h1DA: 	rd_addr = 16'h01D9;      
         12'h1DB: 	rd_addr = 16'h01DA;      
         12'h1DC: 	rd_addr = 16'h01DB;      
         12'h1DD: 	rd_addr = 16'h01DC;      
         12'h1DE: 	rd_addr = 16'h01DD;      
         12'h1DF: 	rd_addr = 16'h01DE;      
         12'h1E0: 	rd_addr = 16'h01DF;      
         12'h1E1:    rd_addr = 16'h01E0;      
         12'h1E2: 	rd_addr = 16'h01E1;      
         12'h1E3: 	rd_addr = 16'h01E2;      
         12'h1E4:    rd_addr = 16'h01E3;   	
         12'h1E5:    rd_addr = 16'h01E4;      
         12'h1E6:  	rd_addr = 16'h01E5;      
         12'h1E7: 	rd_addr = 16'h01E6;      
         12'h1E8: 	rd_addr = 16'h01E7;      
         12'h1E9: 	rd_addr = 16'h01E8;      
         12'h1EA: 	rd_addr = 16'h01E9;      
         12'h1EB: 	rd_addr = 16'h01EA;      
         12'h1EC: 	rd_addr = 16'h01EB;      
         12'h1ED: 	rd_addr = 16'h01EC;      
         12'h1EE: 	rd_addr = 16'h01ED;      
         12'h1EF: 	rd_addr = 16'h01EE;      
         12'h1F0: 	rd_addr = 16'h01EF;      
         12'h1F1: 	rd_addr = 16'h01F0;      
         12'h1F2: 	rd_addr = 16'h01F1;      
         12'h1F3: 	rd_addr = 16'h01F2;      
         12'h1F4: 	rd_addr = 16'h01F3;      
         12'h1F5:    rd_addr = 16'h01F4;      
         12'h1F6:  	rd_addr = 16'h01F5;      
         12'h1F7: 	rd_addr = 16'h01F6;      
         12'h1F8: 	rd_addr = 16'h01F7;      
         12'h1F9: 	rd_addr = 16'h01F8;      
         12'h1FA: 	rd_addr = 16'h01F9;      
         12'h1FB: 	rd_addr = 16'h01FA;      
         12'h1FC: 	rd_addr = 16'h01FB;      
         12'h1FD: 	rd_addr = 16'h01FC;      
         12'h1FE: 	rd_addr = 16'h01FD;      
         12'h1FF: 	rd_addr = 16'h01FE;      
         12'h200:    rd_addr = 16'h01FF;
         12'h201: 	rd_addr = 16'h0200;   
         12'h202: 	rd_addr = 16'h0201;   
         12'h203: 	rd_addr = 16'h0202;   
         12'h204: 	rd_addr = 16'h0203;   
         12'h205: 	rd_addr = 16'h0204;   
         12'h206: 	rd_addr = 16'h0205;   
         12'h207: 	rd_addr = 16'h0206;   
         12'h208: 	rd_addr = 16'h0207;   
         12'h209: 	rd_addr = 16'h0208;   
         12'h20A: 	rd_addr = 16'h0209;   
         12'h20B: 	rd_addr = 16'h020A;   
         12'h20C: 	rd_addr = 16'h020B;   
         12'h20D: 	rd_addr = 16'h020C;   
         12'h20E: 	rd_addr = 16'h020D;   
         12'h20F: 	rd_addr = 16'h020E;   
         12'h210: 	rd_addr = 16'h020F;   
         12'h211: 	rd_addr = 16'h0210;   
         12'h212: 	rd_addr = 16'h0211;   
         12'h213: 	rd_addr = 16'h0212;   
         12'h214: 	rd_addr = 16'h0213;   
         12'h215: 	rd_addr = 16'h0214;   
         12'h216: 	rd_addr = 16'h0215;   
         12'h217: 	rd_addr = 16'h0216;   
         12'h218: 	rd_addr = 16'h0217;   
         12'h219: 	rd_addr = 16'h0218;   
         12'h21A: 	rd_addr = 16'h0219;   
         12'h21B: 	rd_addr = 16'h021A;   
         12'h21C: 	rd_addr = 16'h021B;   
         12'h21D: 	rd_addr = 16'h021C;   
         12'h21E: 	rd_addr = 16'h021D;   
         12'h21F: 	rd_addr = 16'h021E;   
         12'h220: 	rd_addr = 16'h021F;   
         12'h221: 	rd_addr = 16'h0220;   
         12'h222: 	rd_addr = 16'h0221;   
         12'h223: 	rd_addr = 16'h0222;   
         12'h224: 	rd_addr = 16'h0223;   
         12'h225: 	rd_addr = 16'h0224;   
         12'h226: 	rd_addr = 16'h0225;   
         12'h227: 	rd_addr = 16'h0226;   
         12'h228: 	rd_addr = 16'h0227;   
         12'h229: 	rd_addr = 16'h0228;   
         12'h22A: 	rd_addr = 16'h0229;   
         12'h22B: 	rd_addr = 16'h022A;   
         12'h22C: 	rd_addr = 16'h022B;   
         12'h22D: 	rd_addr = 16'h022C;   
         12'h22E: 	rd_addr = 16'h022D;   
         12'h22F: 	rd_addr = 16'h022E;   
         12'h230:    rd_addr = 16'h022F;
         12'h231: 	rd_addr = 16'h0230;   
         12'h232: 	rd_addr = 16'h0231;   
         12'h233: 	rd_addr = 16'h0232;   
         12'h234: 	rd_addr = 16'h0233;   
         12'h235: 	rd_addr = 16'h0234;   
         12'h236: 	rd_addr = 16'h0235;   
         12'h237: 	rd_addr = 16'h0236;   
         12'h238: 	rd_addr = 16'h0237;   
         12'h239: 	rd_addr = 16'h0238;   
         12'h23A: 	rd_addr = 16'h0239;   
         12'h23B: 	rd_addr = 16'h023A;   
         12'h23C: 	rd_addr = 16'h023B;   
         12'h23D: 	rd_addr = 16'h023C;   
         12'h23E: 	rd_addr = 16'h023D;   
         12'h23F: 	rd_addr = 16'h023E;   
         12'h240: 	rd_addr = 16'h023F;   
         12'h241: 	rd_addr = 16'h0240;   
         12'h242: 	rd_addr = 16'h0241;   
         12'h243: 	rd_addr = 16'h0242;   
         12'h244: 	rd_addr = 16'h0243;   
         12'h245: 	rd_addr = 16'h0244;   
         12'h246: 	rd_addr = 16'h0245;   
         12'h247: 	rd_addr = 16'h0246;   
         12'h248: 	rd_addr = 16'h0247;   
         12'h249: 	rd_addr = 16'h0248;   
         12'h24A: 	rd_addr = 16'h0249;   
         12'h24B: 	rd_addr = 16'h024A;   
         12'h24C: 	rd_addr = 16'h024B;   
         12'h24D: 	rd_addr = 16'h024C;   
         12'h24E: 	rd_addr = 16'h024D;   
         12'h24F: 	rd_addr = 16'h024E;   
         12'h250: 	rd_addr = 16'h024F;   
         12'h251: 	rd_addr = 16'h0250;   
         12'h252: 	rd_addr = 16'h0251;   
         12'h253: 	rd_addr = 16'h0252;   
         12'h254: 	rd_addr = 16'h0253;   
         12'h255: 	rd_addr = 16'h0254;   
         12'h256: 	rd_addr = 16'h0255;   
         12'h257: 	rd_addr = 16'h0256;   
         12'h258: 	rd_addr = 16'h0257;   
         12'h259: 	rd_addr = 16'h0258;   
         12'h25A: 	rd_addr = 16'h0259;   
         12'h25B: 	rd_addr = 16'h025A;   
         12'h25C: 	rd_addr = 16'h025B;   
         12'h25D: 	rd_addr = 16'h025C;   
         12'h25E: 	rd_addr = 16'h025D;   
         12'h25F: 	rd_addr = 16'h025E;   
         12'h260: 	rd_addr = 16'h025F;   
         12'h261: 	rd_addr = 16'h0260;   
         12'h262: 	rd_addr = 16'h0261;   
         12'h263:    rd_addr = 16'h0262;  
         12'h264:    rd_addr = 16'h0263;  
         12'h265:    rd_addr = 16'h0264;  
         12'h266:    rd_addr = 16'h0265;  
         12'h267:    rd_addr = 16'h0266;  
         12'h268: 	rd_addr = 16'h0267;      
         12'h269: 	rd_addr = 16'h0268;      
         12'h26A: 	rd_addr = 16'h0269;      
         12'h26B: 	rd_addr = 16'h026A;      
         12'h26C: 	rd_addr = 16'h026B;      
         12'h26D: 	rd_addr = 16'h026C;      
         12'h26E: 	rd_addr = 16'h026D;      
         12'h26F: 	rd_addr = 16'h026E;      
         12'h270:    rd_addr = 16'h026F;   
         12'h271: 	rd_addr = 16'h0270;      
         12'h272: 	rd_addr = 16'h0271;      
         12'h273: 	rd_addr = 16'h0272;      
         12'h274: 	rd_addr = 16'h0273;      
         12'h275: 	rd_addr = 16'h0274;      
         12'h276:    rd_addr = 16'h0275;    
         12'h277:    rd_addr = 16'h0276;    
         12'h278: 	rd_addr = 16'h0277;      
         12'h279: 	rd_addr = 16'h0278;   
         12'h27A:    rd_addr = 16'h0279;       	
         12'h27B:    rd_addr = 16'h027A;    	
         12'h27C:    rd_addr = 16'h027B; 	
         12'h27D: 	rd_addr = 16'h027C;   
         12'h27E: 	rd_addr = 16'h027D;   
         12'h27F: 	rd_addr = 16'h027E;   
         12'h280:    rd_addr = 16'h027F;
         12'h281: 	rd_addr = 16'h0280;   
         12'h282: 	rd_addr = 16'h0281;   
         12'h283: 	rd_addr = 16'h0282;   
         12'h284: 	rd_addr = 16'h0283;   
         12'h285: 	rd_addr = 16'h0284;   
         12'h286:    rd_addr = 16'h0285; 
         12'h287:    rd_addr = 16'h0286; 
         12'h288: 	rd_addr = 16'h0287;   
         12'h289: 	rd_addr = 16'h0288;   
         12'h28A: 	rd_addr = 16'h0289;   
         12'h28B: 	rd_addr = 16'h028A;   
         12'h28C: 	rd_addr = 16'h028B;   
         12'h28D: 	rd_addr = 16'h028C;   
         12'h28E: 	rd_addr = 16'h028D;   
         12'h28F: 	rd_addr = 16'h028E;   
         12'h290:    rd_addr = 16'h028F; 
         12'h291:    rd_addr = 16'h0290;	 
         12'h292: 	rd_addr = 16'h0291;   
         12'h293: 	rd_addr = 16'h0292;   
         12'h294: 	rd_addr = 16'h0293;   
         12'h295: 	rd_addr = 16'h0294;   
         12'h296:    rd_addr = 16'h0295;
         12'h297:    rd_addr = 16'h0296;
         12'h298: 	rd_addr = 16'h0297;
         12'h299: 	rd_addr = 16'h0298;   
         12'h29A: 	rd_addr = 16'h0299;   
         12'h29B:  	rd_addr = 16'h029A;      
         12'h29C: 	rd_addr = 16'h029B;      
         12'h29D: 	rd_addr = 16'h029C;      
         12'h29E: 	rd_addr = 16'h029D;      
         12'h29F: 	rd_addr = 16'h029E;      
         12'h2A0:    rd_addr = 16'h029F;    
         12'h2A1:    rd_addr = 16'h02A0;          	
         12'h2A2:    rd_addr = 16'h02A1; 	
         12'h2A3: 	rd_addr = 16'h02A2;      
         12'h2A4: 	rd_addr = 16'h02A3;      
         12'h2A5: 	rd_addr = 16'h02A4;      
         12'h2A6:    rd_addr = 16'h02A5;    
         12'h2A7:    rd_addr = 16'h02A6;    
         12'h2A8: 	rd_addr = 16'h02A7;      
         12'h2A9: 	rd_addr = 16'h02A8;      
         12'h2AA:    rd_addr = 16'h02A9;	      
         12'h2AB: 	rd_addr = 16'h02AA;      
         12'h2AC: 	rd_addr = 16'h02AB;      
         12'h2AD: 	rd_addr = 16'h02AC;      
         12'h2AE: 	rd_addr = 16'h02AD;      
         12'h2AF: 	rd_addr = 16'h02AE;      
         12'h2B0: 	rd_addr = 16'h02AF;      
         12'h2B1: 	rd_addr = 16'h02B0;      
         12'h2B2: 	rd_addr = 16'h02B1;      
         12'h2B3: 	rd_addr = 16'h02B2;      
         12'h2B4: 	rd_addr = 16'h02B3;      
         12'h2B5:    rd_addr = 16'h02B4;    
         12'h2B6:    rd_addr = 16'h02B5;    
         12'h2B7: 	rd_addr = 16'h02B6;      
         12'h2B8: 	rd_addr = 16'h02B7;      
         12'h2B9: 	rd_addr = 16'h02B8;      
         12'h2BA: 	rd_addr = 16'h02B9;      
         12'h2BB:    rd_addr = 16'h02BA;    	
         12'h2BC:    rd_addr = 16'h02BB;    
         12'h2BD: 	rd_addr = 16'h02BC;      
         12'h2BE: 	rd_addr = 16'h02BD;      
         12'h2BF: 	rd_addr = 16'h02BE;      
         12'h2C0: 	rd_addr = 16'h02BF;      
         12'h2C1: 	rd_addr = 16'h02C0;      
         12'h2C2: 	rd_addr = 16'h02C1;      
         12'h2C3: 	rd_addr = 16'h02C2;      
         12'h2C4: 	rd_addr = 16'h02C3;      
         12'h2C5:    rd_addr = 16'h02C4;    
         12'h2C6:    rd_addr = 16'h02C5;    
         12'h2C7: 	rd_addr = 16'h02C6;      
         12'h2C8: 	rd_addr = 16'h02C7;      
         12'h2C9: 	rd_addr = 16'h02C8;      
         12'h2CA: 	rd_addr = 16'h02C9;      
         12'h2CB: 	rd_addr = 16'h02CA;      
         12'h2CC: 	rd_addr = 16'h02CB;      
         12'h2CD: 	rd_addr = 16'h02CC;      
         12'h2CE: 	rd_addr = 16'h02CD;      
         12'h2CF: 	rd_addr = 16'h02CE;      
         12'h2D0: 	rd_addr = 16'h02CF;      
         12'h2D1: 	rd_addr = 16'h02D0;      
         12'h2D2: 	rd_addr = 16'h02D1;         
         12'h2D3: 	rd_addr = 16'h02D2;      
         12'h2D4: 	rd_addr = 16'h02D3;      
         12'h2D5:    rd_addr = 16'h02D4;    
         12'h2D6:    rd_addr = 16'h02D5;    
         12'h2D7:    rd_addr = 16'h02D6;    	
         12'h2D8: 	rd_addr = 16'h02D7;      
         12'h2D9: 	rd_addr = 16'h02D8;      
         12'h2DA: 	rd_addr = 16'h02D9;      
         12'h2DB: 	rd_addr = 16'h02DA;      
         12'h2DC: 	rd_addr = 16'h02DB;      
         12'h2DD: 	rd_addr = 16'h02DC;      
         12'h2DE: 	rd_addr = 16'h02DD;      
         12'h2DF: 	rd_addr = 16'h02DE;      
         12'h2E0: 	rd_addr = 16'h02DF;      
         12'h2E1:    rd_addr = 16'h02E0;   
         12'h2E2: 	rd_addr = 16'h02E1;      
         12'h2E3: 	rd_addr = 16'h02E2;      
         12'h2E4:    rd_addr = 16'h02E3; 	
         12'h2E5:    rd_addr = 16'h02E4;    
         12'h2E6:    rd_addr = 16'h02E5;    
         12'h2E7: 	rd_addr = 16'h02E6;      
         12'h2E8: 	rd_addr = 16'h02E7;      
         12'h2E9: 	rd_addr = 16'h02E8;      
         12'h2EA: 	rd_addr = 16'h02E9;      
         12'h2EB: 	rd_addr = 16'h02EA;      
         12'h2EC: 	rd_addr = 16'h02EB;      
         12'h2ED: 	rd_addr = 16'h02EC;      
         12'h2EE: 	rd_addr = 16'h02ED;      
         12'h2EF: 	rd_addr = 16'h02EE;      
         12'h2F0: 	rd_addr = 16'h02EF;      
         12'h2F1: 	rd_addr = 16'h02F0;      
         12'h2F2: 	rd_addr = 16'h02F1;      
         12'h2F3: 	rd_addr = 16'h02F2;      
         12'h2F4: 	rd_addr = 16'h02F3;      
         12'h2F5:    rd_addr = 16'h02F4;    
         12'h2F6:    rd_addr = 16'h02F5;    
         12'h2F7: 	rd_addr = 16'h02F6;      
         12'h2F8: 	rd_addr = 16'h02F7;      
         12'h2F9: 	rd_addr = 16'h02F8;      
         12'h2FA:    rd_addr = 16'h02F9;	      
         12'h2FB: 	rd_addr = 16'h02FA;      
         12'h2FC: 	rd_addr = 16'h02FB;      
         12'h2FD: 	rd_addr = 16'h02FC;      
         12'h2FE: 	rd_addr = 16'h02FD;      
         12'h2FF: 	rd_addr = 16'h02FE;      
         12'h300:    rd_addr = 16'h02FF;
         12'h301: 	rd_addr = 16'h0300;   
         12'h302: 	rd_addr = 16'h0301;   
         12'h303: 	rd_addr = 16'h0302;   
         12'h304: 	rd_addr = 16'h0303;   
         12'h305: 	rd_addr = 16'h0304;   
         12'h306: 	rd_addr = 16'h0305;   
         12'h307: 	rd_addr = 16'h0306;   
         12'h308: 	rd_addr = 16'h0307;   
         12'h309: 	rd_addr = 16'h0308;   
         12'h30A: 	rd_addr = 16'h0309;   
         12'h30B: 	rd_addr = 16'h030A;   
         12'h30C: 	rd_addr = 16'h030B;   
         12'h30D: 	rd_addr = 16'h030C;   
         12'h30E: 	rd_addr = 16'h030D;   
         12'h30F: 	rd_addr = 16'h030E;   
         12'h310: 	rd_addr = 16'h030F;   
         12'h311: 	rd_addr = 16'h0310;   
         12'h312: 	rd_addr = 16'h0311;   
         12'h313: 	rd_addr = 16'h0312;   
         12'h314: 	rd_addr = 16'h0313;   
         12'h315: 	rd_addr = 16'h0314;   
         12'h316: 	rd_addr = 16'h0315;   
         12'h317: 	rd_addr = 16'h0316;   
         12'h318: 	rd_addr = 16'h0317;   
         12'h319: 	rd_addr = 16'h0318;   
         12'h31A: 	rd_addr = 16'h0319;   
         12'h31B: 	rd_addr = 16'h031A;   
         12'h31C: 	rd_addr = 16'h031B;   
         12'h31D: 	rd_addr = 16'h031C;   
         12'h31E: 	rd_addr = 16'h031D;   
         12'h31F: 	rd_addr = 16'h031E;   
         12'h320: 	rd_addr = 16'h031F;   
         12'h321: 	rd_addr = 16'h0320;   
         12'h322: 	rd_addr = 16'h0321;   
         12'h323: 	rd_addr = 16'h0322;   
         12'h324: 	rd_addr = 16'h0323;   
         12'h325: 	rd_addr = 16'h0324;   
         12'h326: 	rd_addr = 16'h0325;   
         12'h327: 	rd_addr = 16'h0326;   
         12'h328: 	rd_addr = 16'h0327;   
         12'h329: 	rd_addr = 16'h0328;   
         12'h32A: 	rd_addr = 16'h0329;   
         12'h32B: 	rd_addr = 16'h032A;   
         12'h32C: 	rd_addr = 16'h032B;   
         12'h32D: 	rd_addr = 16'h032C;   
         12'h32E: 	rd_addr = 16'h032D;   
         12'h32F: 	rd_addr = 16'h032E;   
         12'h330:    rd_addr = 16'h032F;
         12'h331: 	rd_addr = 16'h0330;   
         12'h332: 	rd_addr = 16'h0331;   
         12'h333: 	rd_addr = 16'h0332;   
         12'h334: 	rd_addr = 16'h0333;   
         12'h335: 	rd_addr = 16'h0334;   
         12'h336: 	rd_addr = 16'h0335;   
         12'h337: 	rd_addr = 16'h0336;   
         12'h338: 	rd_addr = 16'h0337;   
         12'h339: 	rd_addr = 16'h0338;   
         12'h33A: 	rd_addr = 16'h0339;   
         12'h33B: 	rd_addr = 16'h033A;   
         12'h33C: 	rd_addr = 16'h033B;   
         12'h33D: 	rd_addr = 16'h033C;   
         12'h33E: 	rd_addr = 16'h033D;   
         12'h33F: 	rd_addr = 16'h033E;   
         12'h340: 	rd_addr = 16'h033F;   
         12'h341: 	rd_addr = 16'h0340;   
         12'h342: 	rd_addr = 16'h0341;   
         12'h343: 	rd_addr = 16'h0342;   
         12'h344: 	rd_addr = 16'h0343;   
         12'h345: 	rd_addr = 16'h0344;   
         12'h346: 	rd_addr = 16'h0345;   
         12'h347: 	rd_addr = 16'h0346;   
         12'h348: 	rd_addr = 16'h0347;   
         12'h349: 	rd_addr = 16'h0348;   
         12'h34A: 	rd_addr = 16'h0349;   
         12'h34B: 	rd_addr = 16'h034A;   
         12'h34C: 	rd_addr = 16'h034B;   
         12'h34D: 	rd_addr = 16'h034C;   
         12'h34E: 	rd_addr = 16'h034D;   
         12'h34F: 	rd_addr = 16'h034E;   
         12'h350: 	rd_addr = 16'h034F;   
         12'h351: 	rd_addr = 16'h0350;   
         12'h352: 	rd_addr = 16'h0351;   
         12'h353: 	rd_addr = 16'h0352;   
         12'h354: 	rd_addr = 16'h0353;   
         12'h355: 	rd_addr = 16'h0354;   
         12'h356: 	rd_addr = 16'h0355;   
         12'h357: 	rd_addr = 16'h0356;   
         12'h358: 	rd_addr = 16'h0357;   
         12'h359: 	rd_addr = 16'h0358;   
         12'h35A: 	rd_addr = 16'h0359;   
         12'h35B: 	rd_addr = 16'h035A;   
         12'h35C: 	rd_addr = 16'h035B;   
         12'h35D: 	rd_addr = 16'h035C;   
         12'h35E: 	rd_addr = 16'h035D;   
         12'h35F: 	rd_addr = 16'h035E;   
         12'h360: 	rd_addr = 16'h035F;   
         12'h361: 	rd_addr = 16'h0360;   
         12'h362: 	rd_addr = 16'h0361;   
         12'h363:    rd_addr = 16'h0362;  
         12'h364:    rd_addr = 16'h0363;  
         12'h365:    rd_addr = 16'h0364;  
         12'h366:    rd_addr = 16'h0365;  
         12'h367:    rd_addr = 16'h0366;  
         12'h368: 	rd_addr = 16'h0367;      
         12'h369: 	rd_addr = 16'h0368;      
         12'h36A: 	rd_addr = 16'h0369;      
         12'h36B: 	rd_addr = 16'h036A;      
         12'h36C: 	rd_addr = 16'h036B;      
         12'h36D: 	rd_addr = 16'h036C;      
         12'h36E: 	rd_addr = 16'h036D;      
         12'h36F: 	rd_addr = 16'h036E;      
         12'h370:    rd_addr = 16'h036F;   
         12'h371: 	rd_addr = 16'h0370;      
         12'h372: 	rd_addr = 16'h0371;      
         12'h373: 	rd_addr = 16'h0372;      
         12'h374: 	rd_addr = 16'h0373;      
         12'h375: 	rd_addr = 16'h0374;      
         12'h376:    rd_addr = 16'h0375;    
         12'h377:    rd_addr = 16'h0376;    
         12'h378: 	rd_addr = 16'h0377;      
         12'h379: 	rd_addr = 16'h0378;   
         12'h37A:    rd_addr = 16'h0379;       	
         12'h37B:    rd_addr = 16'h037A;    	
         12'h37C:    rd_addr = 16'h037B; 	
         12'h37D: 	rd_addr = 16'h037C;   
         12'h37E: 	rd_addr = 16'h037D;   
         12'h37F: 	rd_addr = 16'h037E;   
         12'h380:    rd_addr = 16'h037F;
         12'h381: 	rd_addr = 16'h0380;   
         12'h382: 	rd_addr = 16'h0381;   
         12'h383: 	rd_addr = 16'h0382;   
         12'h384: 	rd_addr = 16'h0383;   
         12'h385: 	rd_addr = 16'h0384;   
         12'h386:    rd_addr = 16'h0385; 
         12'h387:    rd_addr = 16'h0386; 
         12'h388: 	rd_addr = 16'h0387;   
         12'h389: 	rd_addr = 16'h0388;   
         12'h38A: 	rd_addr = 16'h0389;   
         12'h38B: 	rd_addr = 16'h038A;   
         12'h38C: 	rd_addr = 16'h038B;   
         12'h38D: 	rd_addr = 16'h038C;   
         12'h38E: 	rd_addr = 16'h038D;   
         12'h38F: 	rd_addr = 16'h038E;   
         12'h390:    rd_addr = 16'h038F; 
         12'h391:    rd_addr = 16'h0390;	 
         12'h392: 	rd_addr = 16'h0391;   
         12'h393: 	rd_addr = 16'h0392;   
         12'h394: 	rd_addr = 16'h0393;   
         12'h395: 	rd_addr = 16'h0394;   
         12'h396:    rd_addr = 16'h0395;
         12'h397:    rd_addr = 16'h0396;
         12'h398: 	rd_addr = 16'h0397;
         12'h399: 	rd_addr = 16'h0398;   
         12'h39A: 	rd_addr = 16'h0399;   
         12'h39B:  	rd_addr = 16'h039A;      
         12'h39C: 	rd_addr = 16'h039B;      
         12'h39D: 	rd_addr = 16'h039C;      
         12'h39E: 	rd_addr = 16'h039D;      
         12'h39F: 	rd_addr = 16'h039E;      
         12'h3A0:    rd_addr = 16'h039F;    
         12'h3A1:    rd_addr = 16'h03A0;          	
         12'h3A2:    rd_addr = 16'h03A1; 	
         12'h3A3: 	rd_addr = 16'h03A2;      
         12'h3A4: 	rd_addr = 16'h03A3;      
         12'h3A5: 	rd_addr = 16'h03A4;      
         12'h3A6:    rd_addr = 16'h03A5;    
         12'h3A7:    rd_addr = 16'h03A6;    
         12'h3A8: 	rd_addr = 16'h03A7;      
         12'h3A9: 	rd_addr = 16'h03A8;      
         12'h3AA:    rd_addr = 16'h03A9;	      
         12'h3AB: 	rd_addr = 16'h03AA;      
         12'h3AC: 	rd_addr = 16'h03AB;      
         12'h3AD: 	rd_addr = 16'h03AC;      
         12'h3AE: 	rd_addr = 16'h03AD;      
         12'h3AF: 	rd_addr = 16'h03AE;      
         12'h3B0: 	rd_addr = 16'h03AF;      
         12'h3B1: 	rd_addr = 16'h03B0;      
         12'h3B2: 	rd_addr = 16'h03B1;      
         12'h3B3: 	rd_addr = 16'h03B2;      
         12'h3B4: 	rd_addr = 16'h03B3;      
         12'h3B5:    rd_addr = 16'h03B4;    
         12'h3B6:    rd_addr = 16'h03B5;    
         12'h3B7: 	rd_addr = 16'h03B6;      
         12'h3B8: 	rd_addr = 16'h03B7;      
         12'h3B9: 	rd_addr = 16'h03B8;      
         12'h3BA: 	rd_addr = 16'h03B9;      
         12'h3BB:    rd_addr = 16'h03BA;    	
         12'h3BC:    rd_addr = 16'h03BB;    
         12'h3BD: 	rd_addr = 16'h03BC;      
         12'h3BE: 	rd_addr = 16'h03BD;      
         12'h3BF: 	rd_addr = 16'h03BE;      
         12'h3C0: 	rd_addr = 16'h03BF;      
         12'h3C1: 	rd_addr = 16'h03C0;      
         12'h3C2: 	rd_addr = 16'h03C1;      
         12'h3C3: 	rd_addr = 16'h03C2;      
         12'h3C4: 	rd_addr = 16'h03C3;      
         12'h3C5:    rd_addr = 16'h03C4;    
         12'h3C6:    rd_addr = 16'h03C5;    
         12'h3C7: 	rd_addr = 16'h03C6;      
         12'h3C8: 	rd_addr = 16'h03C7;      
         12'h3C9: 	rd_addr = 16'h03C8;      
         12'h3CA: 	rd_addr = 16'h03C9;      
         12'h3CB: 	rd_addr = 16'h03CA;      
         12'h3CC: 	rd_addr = 16'h03CB;      
         12'h3CD: 	rd_addr = 16'h03CC;      
         12'h3CE: 	rd_addr = 16'h03CD;      
         12'h3CF: 	rd_addr = 16'h03CE;      
         12'h3D0: 	rd_addr = 16'h03CF;      
         12'h3D1: 	rd_addr = 16'h03D0;      
         12'h3D2: 	rd_addr = 16'h03D1;         
         12'h3D3: 	rd_addr = 16'h03D2;      
         12'h3D4: 	rd_addr = 16'h03D3;      
         12'h3D5:    rd_addr = 16'h03D4;    
         12'h3D6:    rd_addr = 16'h03D5;    
         12'h3D7:    rd_addr = 16'h03D6;    	
         12'h3D8: 	rd_addr = 16'h03D7;      
         12'h3D9: 	rd_addr = 16'h03D8;      
         12'h3DA: 	rd_addr = 16'h03D9;      
         12'h3DB: 	rd_addr = 16'h03DA;      
         12'h3DC: 	rd_addr = 16'h03DB;      
         12'h3DD: 	rd_addr = 16'h03DC;      
         12'h3DE: 	rd_addr = 16'h03DD;      
         12'h3DF: 	rd_addr = 16'h03DE;      
         12'h3E0: 	rd_addr = 16'h03DF;      
         12'h3E1:    rd_addr = 16'h03E0;   
         12'h3E2: 	rd_addr = 16'h03E1;      
         12'h3E3: 	rd_addr = 16'h03E2;      
         12'h3E4:    rd_addr = 16'h03E3; 	
         12'h3E5:    rd_addr = 16'h03E4;    
         12'h3E6:    rd_addr = 16'h03E5;    
         12'h3E7: 	rd_addr = 16'h03E6;      
         12'h3E8: 	rd_addr = 16'h03E7;      
         12'h3E9: 	rd_addr = 16'h03E8;      
         12'h3EA: 	rd_addr = 16'h03E9;      
         12'h3EB: 	rd_addr = 16'h03EA;      
         12'h3EC: 	rd_addr = 16'h03EB;      
         12'h3ED: 	rd_addr = 16'h03EC;      
         12'h3EE: 	rd_addr = 16'h03ED;      
         12'h3EF: 	rd_addr = 16'h03EE;      
         12'h3F0: 	rd_addr = 16'h03EF;      
         12'h3F1: 	rd_addr = 16'h03F0;      
         12'h3F2: 	rd_addr = 16'h03F1;      
         12'h3F3: 	rd_addr = 16'h03F2;      
         12'h3F4: 	rd_addr = 16'h03F3;      
         12'h3F5:    rd_addr = 16'h03F4;    
         12'h3F6:    rd_addr = 16'h03F5;    
         12'h3F7: 	rd_addr = 16'h03F6;      
         12'h3F8: 	rd_addr = 16'h03F7;      
         12'h3F9: 	rd_addr = 16'h03F8;      
         12'h3FA:    rd_addr = 16'h03F9;	      
         12'h3FB: 	rd_addr = 16'h03FA;      
         12'h3FC: 	rd_addr = 16'h03FB;      
         12'h3FD: 	rd_addr = 16'h03FC;      
         12'h3FE: 	rd_addr = 16'h03FD;      
         12'h3FF: 	rd_addr = 16'h03FE;      
         //12'h400:    rd_addr = 16'h03FF;      
         12'h400:    rd_addr = 16'h0123;
			default:	   rd_addr = 16'h0023;
      endcase
					
endmodule
